module OurAdder ( // This is a template. 
// You can modify the input-output declerations(width etc.) without changing the names.
    input[3:0] a, // input A
    input[3:0] b, // input B
    output[3:0] sum // sum output
);

assign sum = a + b;

endmodule
